    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine #�^\     �    bplist00�3A�mQ�*
                            bplist00�_�https://doc-0s-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/1j4ikks06g5p5euo4vun1baha9hvrm93/1549699200000/03251620456578107196/03251620456578107196/1uZNCRDs0EUN2oVGBK0JGjLd41c87-op0?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea323;Safari;9BE98101-3ECF-41B6-90B1-8E06E048B90C 