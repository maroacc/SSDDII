    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine :�^\    8 z"    bplist00�3A�m]I;m
                            bplist00�_�https://doc-08-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/215vao6j0v5h7d256l874ao868vodgnk/1549699200000/03251620456578107196/03251620456578107196/1ROqpehzilrOAj32CS52htzWiMz3pQZQW?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea33a;Safari;9BAA4E60-87F1-4DF1-8AA8-3FD6B61F3D00 