    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine .�^\    �M�"    bplist00�3A�mWH%�
                            bplist00�_�https://doc-0c-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/ieio06ulj7qn7vn4f6nqf2sn633m9tvf/1549699200000/03251620456578107196/03251620456578107196/1dBxppAZIFhE98MaO5KXOjyLxXlXrGcqg?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea32e;Safari;1E7A253C-10B5-446B-B65E-42639D88A35E 