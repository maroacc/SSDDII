    Mac OS X            	   2  ,     ^                                      ATTR      ^  $  :                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  �  %com.apple.metadata:kMDItemWhereFroms   "   <  com.apple.quarantine �^\     �    bplist00�3A�mJ�l�
                            bplist00�_5https://doc-00-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/anem8vlaill1ajp2ugqtmts6mjv35bkl/1549699200000/03251620456578107196/03251620456578107196/1yO3Intyc47NQqxOa_TIiaBFb484G5V6e?e=download&nonce=po0mrgapu1qec&user=03251620456578107196&hash=4j1drdjkhhddg89f4qplepba4k56njso_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP  D                           �q/0083;5c5ea315;Safari;90900B83-B35E-4426-8002-1EE426BD6743 