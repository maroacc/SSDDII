    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine %�^\    ?Z    bplist00�3A�mR��4
                            bplist00�_�https://doc-0c-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/lg4lq6bced23ekti0ui720b84fjakq36/1549699200000/03251620456578107196/03251620456578107196/1zeX0rDpGEU0WeqJesVs2wh8bOPa3K2Aa?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea325;Safari;A6FE7BA1-0053-4B0F-899F-CF790F583D80 