    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine +�^\    =M&    bplist00�3A�mU�i�
                            bplist00�_�https://doc-00-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/a2m83bt7scrleqlia7u41ob1i68ufvea/1549699200000/03251620456578107196/03251620456578107196/1qwY0yUW6_6X72WDDwiHVQ55Wr2sUADik?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea32b;Safari;5836EC36-5D77-4163-ABF7-22B5E5E42476 