    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine )�^\    �r�    bplist00�3A�mT�'�
                            bplist00�_�https://doc-14-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/lebld2nct9fi4l4h4ancc65cjj3m1dbr/1549699200000/03251620456578107196/03251620456578107196/1YxeK4izmvbPcWrJYf9z3Qaa73Lt0kCxL?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea329;Safari;13C68CB5-A779-4002-BFB1-4C0E52E058D8 