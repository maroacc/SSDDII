    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine 7�^\    x��+    bplist00�3A�m[�\>
                            bplist00�_�https://doc-0s-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/el5gnk8bvv4f99j9i6u92e5ktmgnje9n/1549699200000/03251620456578107196/03251620456578107196/1GncDqSg72wQlRJpDhDdQIF6Ssx3z6fQe?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea337;Safari;2B43E7F6-B085-4F12-B6C9-67B36D88891A 