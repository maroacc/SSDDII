    Mac OS X            	   2  �     	                                      ATTR      	  $  �                 $     com.apple.lastuseddate#PS      4   5  )com.apple.metadata:kMDItemDownloadedDate   i  d  %com.apple.metadata:kMDItemWhereFroms   �   <  com.apple.quarantine '�^\    . q    bplist00�3A�mS��
                            bplist00�_�https://doc-0g-bs-docs.googleusercontent.com/docs/securesc/eicg8f771et6jhnt799i37dj9akk4jgb/c6ifrlt4sgieleiqn6mkq31alrqgfj8q/1549699200000/03251620456578107196/03251620456578107196/1Sf_foAEXf8-k9x2AC_GaavQ2_IUFsBWw?e=download_Lhttps://drive.google.com/drive/u/0/folders/1Oxp2RgudZHJvRuAY60eoPttjmdPOQXnP   �                           >q/0083;5c5ea327;Safari;0D4D899A-80EB-4F76-AB79-5EF4007D734C 